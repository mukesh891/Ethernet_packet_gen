class eth_master_sqr extends uvm_sequencer#(eth_seq_item);
  `uvm_component_utils(eth_master_sqr)
  //`NEW_COMP
 function new(string name="", uvm_component parent=null); 
		super.new(name,parent);  
  

  endfunction
     

  
endclass